`timescale 1ns / 1ps

// Mod�l �smi: pulp_clock_gating
// Bu isim, �a��ran dosyadaki (clock_divider) isimle B�REB�R AYNI olmal�d�r.
module pulp_clock_gating (
    input  logic clk_i,
    input  logic en_i,
    input  logic test_en_i,
    output logic clk_o
);

    logic clk_en;

    // -------------------------------------------------------------
    // Latch Tabanl� Clock Gating (Glitch-Free)
    // -------------------------------------------------------------
    // Clock High iken enable de�i�irse ��k��ta "i�ne" (glitch) olu�ur.
    // Latch kullanarak enable sinyalini Clock Low iken g�ncelliyoruz.
    // B�ylece Clock High oldu�unda enable sinyali �oktan sabitlenmi� olur.
    
    always_latch begin
        if (clk_i == 1'b0) begin
            clk_en <= en_i | test_en_i;
        end
    end

    // Saati ge�ir (1) veya kes (0)
    assign clk_o = clk_i & clk_en;

endmodule