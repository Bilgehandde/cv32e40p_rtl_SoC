`timescale 1ns / 1ps

// ========================================================================
// 1. PULP CLOCK MUX 2 (Saat Se�ici)
// ========================================================================
// �ki saat kayna�� aras�nda se�im yapar.
module pulp_clock_mux2 (
    input  logic clk0_i, // Se�im 0
    input  logic clk1_i, // Se�im 1
    input  logic sel_i,  // Se�ici Sinyal
    output logic clk_o   // ��k�� Saati
);
    // Sim�lasyon i�in basit MUX davran���:
    assign clk_o = (sel_i) ? clk1_i : clk0_i;

endmodule

// ========================================================================
// 2. PULP CLOCK XOR 2 (Saat Kar��t�r�c�)
// ========================================================================
// �ki saati XOR i�lemine sokar.
module pulp_clock_xor2 (
    input  logic clk0_i,
    input  logic clk1_i,
    output logic clk_o
);
    assign clk_o = clk0_i ^ clk1_i;

endmodule

// ========================================================================
// 3. PULP CLOCK INVERTER (Saat Tersleyici)
// ========================================================================
// Saatin faz�n� ters �evirir (180 derece).
module pulp_clock_inverter (
    input  logic clk_i,
    output logic clk_o
);
    assign clk_o = ~clk_i;

endmodule